module main

import v.builder.llvmbuilder

fn main() {
	llvmbuilder.start()
}
